<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,121.8,-61.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_INVERTER</type>
<position>14.5,-7.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_INVERTER</type>
<position>15,-33</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>4,-7.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>4,-18</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>4.5,-28.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND3</type>
<position>26.5,-14</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND3</type>
<position>27,-22</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>35,-14</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>35.5,-22</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-7.5,11.5,-7.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-16,23.5,-16</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>17.5 3</intersection>
<intersection>23 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17.5,-16,17.5,-7.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-16 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>23,-24,23,-16</points>
<intersection>-24 5</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23,-24,24,-24</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>23 4</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-22,14.5,-12</points>
<intersection>-22 3</intersection>
<intersection>-18 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-12,23.5,-12</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-18,14.5,-18</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-22,24,-22</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-33,21,-20</points>
<intersection>-33 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-20,24,-20</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-33,21,-33</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-22,34.5,-22</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-14,34,-14</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-28.5,14.5,-14</points>
<intersection>-28.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-14,23.5,-14</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-28.5,14.5,-28.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>11.5 3</intersection>
<intersection>14.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>11.5,-33,11.5,-28.5</points>
<intersection>-33 4</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11.5,-33,12,-33</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>11.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 9></circuit>