<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,121.8,-61.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>3,-3</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>3,-8</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>3,-13.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND3</type>
<position>21.5,-3.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>21.5,-10.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND3</type>
<position>21.5,-17.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND3</type>
<position>21.5,-24</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND3</type>
<position>21.5,-31</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND3</type>
<position>21.5,-38</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND3</type>
<position>21.5,-45</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>BA_NAND3</type>
<position>21.5,-52.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>14.5,-47</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>14.5,-15.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>14.5,-19.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>38.5,-23.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-3,11.5,-1.5</points>
<intersection>-3 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-1.5,18.5,-1.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-3,11.5,-3</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>11,-50.5,11,-1.5</points>
<intersection>-50.5 10</intersection>
<intersection>-43 11</intersection>
<intersection>-36 12</intersection>
<intersection>-29 13</intersection>
<intersection>-22 14</intersection>
<intersection>-15.5 4</intersection>
<intersection>-8.5 15</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11,-15.5,12.5,-15.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>11,-50.5,18.5,-50.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>11,-43,18.5,-43</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>11,-36,18.5,-36</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>11,-29,18.5,-29</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>11,-22,18.5,-22</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>11,-8.5,18.5,-8.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-15.5,18.5,-15.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-19.5,18.5,-19.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-47,18.5,-47</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-8,11.5,-3.5</points>
<intersection>-8 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-8,11.5,-8</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-3.5,18.5,-3.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-52.5,17,-3.5</points>
<intersection>-52.5 10</intersection>
<intersection>-45 11</intersection>
<intersection>-38 12</intersection>
<intersection>-31 13</intersection>
<intersection>-24 14</intersection>
<intersection>-17.5 15</intersection>
<intersection>-10.5 16</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>17,-52.5,18.5,-52.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>17,-45,18.5,-45</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>17,-38,18.5,-38</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>17,-31,18.5,-31</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>17,-24,18.5,-24</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>17,-17.5,18.5,-17.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>17,-10.5,18.5,-10.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-19.5,11.5,-5.5</points>
<intersection>-19.5 4</intersection>
<intersection>-13.5 1</intersection>
<intersection>-12.5 3</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-13.5,11.5,-13.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-5.5,18.5,-5.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11.5,-12.5,18.5,-12.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>11.5,-19.5,18.5,-19.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection>
<intersection>18.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>18.5,-54.5,18.5,-19.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-47 8</intersection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>12.5,-47,18.5,-47</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>18.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-23.5,31,-3.5</points>
<intersection>-23.5 1</intersection>
<intersection>-17.5 4</intersection>
<intersection>-10.5 3</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-23.5,37.5,-23.5</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-3.5,31,-3.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-10.5,31,-10.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-17.5,31,-17.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>24.5 5</intersection>
<intersection>31 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>24.5,-52.5,24.5,-17.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-17.5 4</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,121.8,-61.5</PageViewport></page 9></circuit>